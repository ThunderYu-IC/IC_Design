module hw_1_4 (
    input       [15:0]temp_code,
    output  reg  [7:0]bcd_code
);

always@(temp_code)
begin
    case(temp_code)
        16'b0000_0000_0000_0000: bcd_code = 8'b0000_0000;
        16'b0000_0000_0000_0001: bcd_code = 8'b0000_0001;
        16'b0000_0000_0000_0011: bcd_code = 8'b0000_0010;
        16'b0000_0000_0000_0111: bcd_code = 8'b0000_0011;//3

        16'b0000_0000_0000_1111: bcd_code = 8'b0000_0100;
        16'b0000_0000_0001_1111: bcd_code = 8'b0000_0101;
        16'b0000_0000_0011_1111: bcd_code = 8'b0000_0110;
        16'b0000_0000_0111_1111: bcd_code = 8'b0000_0111;//7

        16'b0000_0000_1111_1111: bcd_code = 8'b0000_1000;
        16'b0000_0001_1111_1111: bcd_code = 8'b0000_1001;
        16'b0000_0011_1111_1111: bcd_code = 8'b0001_0000;
        16'b0000_0111_1111_1111: bcd_code = 8'b0001_0001;//11

        16'b0000_1111_1111_1111: bcd_code = 8'b0001_0010;
        16'b0001_1111_1111_1111: bcd_code = 8'b0001_0011;
        16'b0011_1111_1111_1111: bcd_code = 8'b0001_0100;
        16'b0111_1111_1111_1111: bcd_code = 8'b0001_0101;//15

        16'b1111_1111_1111_1111: bcd_code = 8'b0001_0110;//16
        default: bcd_code = 8'b1111_1111;
    endcase
end    
endmodule

module hw_1_4_2 (
    input       [15:0]I,
    output       [7:0]O
);
    assign O[4] = I[9];
    assign O[3] = ~I[9]&I[7];
    assign O[2] = ( ~I[7]&I[3] | I[13] );
    assign O[1] = ( (~I[3]&I[1]) | (~I[7]&I[5]) | ~(I[13]&I[11]) | I[16] );
    assign O[0] = ( (~I[15]&I[14]) | (~I[13]&I[12]) | (~I[11]&I[10]) | (~I[9]&I[8])
                  | (~I[7]&I[6]) | (~I[5]&I[4]) | (~I[3]&I[2]) | (~I[1]&I[0]) );
endmodule